`timescale 1ns/1ns

module lu3(a, b, op, y);
	input  [7:0] a, b;
	input  [1:0] op;
	output [7:0] y;
	wire   [7:0] w0, w1, w2, w3;
	wire   [3:0] c;
	/* write answer below */
	
	/* write answer above */
endmodule
