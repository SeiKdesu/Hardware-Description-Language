`timescale 1ns/1ns

module stopwatch (clk, rst, sw1, sw2, sw3, dsp);
	input        clk, rst, sw1, sw2, sw3;
	output [7:0] dsp;
	wire ci, ld, clr;

	/* write answer below */

	/* write answer above */

endmodule	
