`timescale 1ns/1ns

module lu2(a, b, op, y);
	input  [7:0] a, b;
	input  [1:0] op;
	output [7:0] y;
	wire   [7:0] w0, w1, w2, w3;
	/* write answer below */
	
	/* write answer above */
endmodule
